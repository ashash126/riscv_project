

`include "defines.v"

// 将指令向译码模块传递
module if_id(

    input wire clk,
    input wire rst,

    input wire[`InstBus] inst_i,            // 指令内容 从指令存储器传入
    input wire[`InstAddrBus] inst_addr_i,   // 指令地址 

    //input wire[`Hold_Flag_Bus] hold_flag_i, // 流水线暂停标志

    input wire rst_if_id_i,             // 复位流水线寄存器信号 

    //input wire[`INT_BUS] int_flag_i,        // 外设中断输入信号
    //output wire[`INT_BUS] int_flag_o,

    output wire[`InstBus] inst_o,           // 指令内容
    output wire[`InstAddrBus] inst_addr_o   // 指令地址

    
    );

    wire[`InstBus] inst;
    gen_pipe_dff #(32) inst_ff(clk, rst, rst_if_id_i, `INST_NOP, inst_i, inst);// 1
    assign inst_o = inst;

    wire[`InstAddrBus] inst_addr;
    gen_pipe_dff #(32) inst_addr_ff(clk, rst, rst_if_id_i, `ZeroWord, inst_addr_i, inst_addr); //0
    assign inst_addr_o = inst_addr;

    //wire[`INT_BUS] int_flag;
    //gen_pipe_dff #(8) int_ff(clk, rst, hold_en, `INT_NONE, int_flag_i, int_flag);
    //assign int_flag_o = int_flag;

endmodule
